LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RAM_32x4_1Port IS
	PORT
	(
		ADDRESS			:	IN		STD_LOGIC_VECTOR	(4 DOWNTO 0);
		DATA_IN			:	IN		STD_LOGIC_VECTOR	(3 DOWNTO 0);
		WRITE_ENABLE	:	IN		STD_LOGIC;
		CLOCK				:	IN		STD_LOGIC;
		DATA_OUT			:	OUT	STD_LOGIC_VECTOR	(3 DOWNTO 0)
	);
END RAM_32x4_1Port;

ARCHITECTURE RAM_32x4 OF RAM_32x4_1Port IS

	TYPE RAM_ARRAY IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL RAM : RAM_ARRAY :=
		(
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0",
			X"0",X"0",X"0",X"0"
		); 

BEGIN

	RAM_1Port : PROCESS(CLOCK)
	BEGIN
		IF(RISING_EDGE(CLOCK)) THEN
			IF(WRITE_ENABLE='1') THEN
				RAM(TO_INTEGER(UNSIGNED(ADDRESS))) <= DATA_IN;
			END IF;
		END IF;
	END PROCESS RAM_1Port;
	
	DATA_OUT <= RAM(TO_INTEGER(UNSIGNED(ADDRESS)));

END RAM_32x4;